`timescale 1ns / 1ps
module wb(
    );


endmodule
